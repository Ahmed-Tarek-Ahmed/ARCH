LIBRARY IEEE;
USE IEEE.std_logic_1164.all;

Entity processor IS 
port(
);
END ENTITY;

Architecture p1 OF processor IS

begin

END Architecture;